package torrence_types;
    typedef int unsigned uint32_t;
    typedef byte unsigned uint8_t;
endpackage
