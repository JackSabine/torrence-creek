typedef struct packed {
    bit is_hit;
    uint32_t req_word;
} cache_response_t;
