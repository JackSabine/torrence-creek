interface reset_if (
    input bit clk
);
    logic reset;
endinterface
