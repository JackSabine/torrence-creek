`include "cache_base_test.sv"
`include "icache_basic_test.sv"
`include "dcache_basic_test.sv"
`include "l1_basic_test.sv"
`include "l1_thrashing_test.sv"
